library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package data_types is
  subtype data_word is signed ( 15 downto  0);
end data_types;

package body data_types is

end data_types;
